module name
#(
    parameter DATA_WIDTH = 32
)
(
    // Inputs
        // Secuential control
            input logic clk,
            input logic async_rst_n,
            input logic sync_rst_n,
            input logic flush,
        // Handshake
        // Data
    // Outputs
        // Handshake
        // Data
);
    import rv32i_types_pkg::*;

endmodule